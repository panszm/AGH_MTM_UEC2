`timescale 1ns / 1ps

module game_board_select
    (   
        input logic clk,
        input logic rst,
        input logic[2:0] board_size,
        input logic[2:0] lvl,
        input logic[1:0] seed,
        output logic[5:0] selected_board [15:0][15:0],
        output logic[5:0] selected_board_complete [15:0][15:0]
    );

    logic [7:0] selection;
    logic[5:0] selected_board_nxt [15:0][15:0];
    logic[5:0] selected_board_complete_nxt [15:0][15:0];
    assign selection = (board_size<<5) + (lvl<<2)+ seed;

    always_ff @(posedge clk) begin
        if(rst) begin
            selected_board <= '{default:0}; 
            selected_board_complete <= '{default:0}; 
        end else begin
            selected_board <= selected_board_nxt;
            selected_board_complete <= selected_board_complete_nxt;
        end
    end

    always_comb begin
case (selection)
            8'b010_001_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000110}
};
                end
            8'b010_001_01: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000100},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000111}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000100},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000111}
};


                end
            8'b010_001_10: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000000, 6'b000111}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001000, 6'b000111}
};


                end
            8'b010_010_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000000, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001000, 6'b000110}
};
                end
            8'b010_010_01: 
                begin
                   selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000100},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000110}
};
                end
            8'b010_010_10: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000000, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000010, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000110}
};
                end
            8'b010_011_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000000, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000000, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000110, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000010, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000110}
};
                end
            8'b010_011_01: 
                begin
                   selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b000000, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b001001, 6'b000111}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000010, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001000, 6'b000011, 6'b000101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000100, 6'b000011, 6'b001001, 6'b000111}
};
                end
            8'b010_011_10: 
                begin
                   selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000000, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000111, 6'b000100, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001001, 6'b000011, 6'b000100},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b001001, 6'b000110}
};
                end
            8'b011_001_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000100}
};
                end
            8'b011_001_01: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b000000, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001000, 6'b000101}
};
                end
            8'b011_001_10: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000000, 6'b001001, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000110, 6'b001001, 6'b000101}
};
                end
            8'b011_010_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b000000, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001000, 6'b000100}
};
                end
            8'b011_010_01: 
                begin
                   selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b000000, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b000000, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001110, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001100, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000101}
};
                end
            8'b011_010_10: 
                begin
                   selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b000000, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001000, 6'b000101}
};
                end
            8'b011_011_00: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b000000, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b000000, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000000}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010000, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001100, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000100}
};
                end
            8'b011_011_01: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b000000, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010010},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000110},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010001, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010011, 6'b001111, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001000, 6'b000101}
};
                end
            8'b011_011_10: 
                begin
                    selected_board_nxt ='{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000101}
};
                    selected_board_complete_nxt = '{
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000101, 6'b000011, 6'b000111, 6'b001011, 6'b001001, 6'b001101, 6'b001111, 6'b010001, 6'b010011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001001, 6'b001011, 6'b001101, 6'b001111, 6'b010001, 6'b010011, 6'b000101, 6'b000011, 6'b000111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001111, 6'b010001, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b001001, 6'b001011, 6'b001101},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000111, 6'b001101, 6'b001001, 6'b010011, 6'b000011, 6'b010001, 6'b001011, 6'b000101, 6'b001111},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000011, 6'b000101, 6'b001111, 6'b001001, 6'b001011, 6'b000111, 6'b001101, 6'b010011, 6'b010001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b001111, 6'b000011, 6'b000111, 6'b001001},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b001101, 6'b000111, 6'b000011, 6'b000101, 6'b010011, 6'b001001, 6'b010001, 6'b001111, 6'b001011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010000, 6'b001001, 6'b000101, 6'b000111, 6'b001111, 6'b001011, 6'b010011, 6'b001101, 6'b000011},
    '{6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b000000, 6'b010010, 6'b001110, 6'b001011, 6'b010001, 6'b001101, 6'b000011, 6'b000111, 6'b001001, 6'b000101}
};
                end
            8'b100_001_00: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b000000 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010100 }};

                end
            8'b100_001_01: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b000000 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010000 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_001_10: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b000000 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100000 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_010_00: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b000000 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b000000, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100000 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010000, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_010_01: 
                begin
                    selected_board_nxt ='{
'{6'b000000, 6'b000000, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001000, 6'b000010, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_010_10: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b000000, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b000000, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011010, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010000, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_011_00: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b000000, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b000000, 6'b001111, 6'b000000, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010010, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011100, 6'b001111, 6'b011000, 6'b001011, 6'b010101 }};

                end
            8'b100_011_01: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b000000 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b000000 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b000000 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001010 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011100 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010000 },
'{6'b010001, 6'b011111, 6'b001001, 6'b000011, 6'b010011, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            8'b100_011_10: 
                begin
                    selected_board_nxt ='{
'{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b000000, 6'b000000, 6'b000000, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                    selected_board_complete_nxt = '{
    '{6'b001001, 6'b000011, 6'b000101, 6'b000111, 6'b001101, 6'b011111, 6'b001111, 6'b011101, 6'b100001, 6'b011011, 6'b010001, 6'b011001, 6'b010111, 6'b010101, 6'b010011, 6'b001011 },
'{6'b010111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001001, 6'b011001, 6'b001011, 6'b011101, 6'b010011, 6'b000011, 6'b000111, 6'b000101, 6'b011111, 6'b001111, 6'b001101 },
'{6'b011111, 6'b001111, 6'b001011, 6'b011001, 6'b000111, 6'b000011, 6'b000101, 6'b001111, 6'b010101, 6'b010111, 6'b001001, 6'b001101, 6'b100001, 6'b010001, 6'b011011, 6'b011101 },
'{6'b011101, 6'b001101, 6'b001111, 6'b010001, 6'b010111, 6'b011011, 6'b100001, 6'b010101, 6'b011111, 6'b001111, 6'b001011, 6'b000101, 6'b000011, 6'b001001, 6'b011001, 6'b000111 },
'{6'b000011, 6'b000101, 6'b010111, 6'b001001, 6'b011001, 6'b010101, 6'b011111, 6'b000111, 6'b010001, 6'b100001, 6'b011101, 6'b001011, 6'b011011, 6'b001111, 6'b001101, 6'b010011 },
'{6'b001101, 6'b011101, 6'b010001, 6'b010101, 6'b001111, 6'b000101, 6'b001001, 6'b011011, 6'b001111, 6'b011001, 6'b000111, 6'b010111, 6'b001011, 6'b100001, 6'b000011, 6'b011111 },
'{6'b001111, 6'b010011, 6'b011011, 6'b001011, 6'b011101, 6'b100001, 6'b010111, 6'b000011, 6'b001101, 6'b010101, 6'b011111, 6'b001001, 6'b011001, 6'b000111, 6'b001101, 6'b000101 },
'{6'b000111, 6'b100001, 6'b011001, 6'b011111, 6'b001011, 6'b010011, 6'b010001, 6'b001101, 6'b000101, 6'b000011, 6'b011011, 6'b001111, 6'b010101, 6'b011101, 6'b001001, 6'b010111 },
'{6'b011011, 6'b001011, 6'b011111, 6'b011101, 6'b001001, 6'b001101, 6'b010101, 6'b010111, 6'b000111, 6'b000101, 6'b011001, 6'b000011, 6'b010001, 6'b010011, 6'b100001, 6'b001111 },
'{6'b011001, 6'b001001, 6'b001111, 6'b001101, 6'b000011, 6'b011101, 6'b010011, 6'b011111, 6'b001011, 6'b010001, 6'b100001, 6'b010101, 6'b000111, 6'b010111, 6'b000101, 6'b011011 },
'{6'b010011, 6'b010001, 6'b000011, 6'b010111, 6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b001111, 6'b011101, 6'b001101, 6'b011011, 6'b011111, 6'b001011, 6'b010101, 6'b001001 },
'{6'b000101, 6'b000111, 6'b010101, 6'b100001, 6'b011011, 6'b010001, 6'b001011, 6'b001111, 6'b001001, 6'b011111, 6'b010111, 6'b010011, 6'b001101, 6'b000011, 6'b011101, 6'b011001 },
'{6'b001011, 6'b010111, 6'b001101, 6'b010011, 6'b011111, 6'b001111, 6'b011011, 6'b010001, 6'b011001, 6'b001001, 6'b010101, 6'b100001, 6'b011101, 6'b000101, 6'b000111, 6'b000011 },
'{6'b010101, 6'b011011, 6'b011101, 6'b001111, 6'b000101, 6'b000111, 6'b000011, 6'b011001, 6'b010111, 6'b001011, 6'b010011, 6'b010001, 6'b001001, 6'b011101, 6'b011111, 6'b100001 },
'{6'b100001, 6'b011001, 6'b000111, 6'b000101, 6'b010101, 6'b001011, 6'b011101, 6'b001001, 6'b000011, 6'b001101, 6'b001111, 6'b011111, 6'b010011, 6'b011011, 6'b010111, 6'b010001 },
'{6'b010001, 6'b011111, 6'b001000, 6'b000010, 6'b010010, 6'b010111, 6'b001101, 6'b100001, 6'b011011, 6'b000111, 6'b000101, 6'b011101, 6'b001111, 6'b011001, 6'b001011, 6'b010101 }};

                end
            default: 
                begin
                    selected_board_nxt = '{default:0}; 

                    selected_board_complete_nxt = '{default:0};
                end
        endcase
    end

endmodule
