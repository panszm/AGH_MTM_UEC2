`timescale 1ns / 1ps
// ROM with synchonous read (inferring Block RAM)
// character ROM
module font_rom_numerical
    (
        input  wire        clk,
        input  wire [10:0] addr,            // {char_code[6:0], char_line[3:0]}
        output reg  [7:0]  char_line_pixels // pixels of the character line
    );

    // signal declaration
    reg [7:0] data;

    // body
    always @(posedge clk)
        char_line_pixels <= data;

    always @*
        case (addr)
            //code x00
            11'h000: data = 8'b00000000; //
            11'h001: data = 8'b00000000; //
            11'h002: data = 8'b00000000; //
            11'h003: data = 8'b00000000; //
            11'h004: data = 8'b00000000; //
            11'h005: data = 8'b00000000; //
            11'h006: data = 8'b00000000; //
            11'h007: data = 8'b00000000; //
            11'h008: data = 8'b00000000; //
            11'h009: data = 8'b00000000; //
            11'h00a: data = 8'b00000000; //
            11'h00b: data = 8'b00000000; //
            11'h00c: data = 8'b00000000; //
            11'h00d: data = 8'b00000000; //
            11'h00e: data = 8'b00000000; //
            11'h00f: data = 8'b00000000; //
            //code x01
            11'h010: data = 8'b00000000; //
            11'h011: data = 8'b00000000; //
            11'h012: data = 8'b01111100; //  *****
            11'h013: data = 8'b11000110; // **   **
            11'h014: data = 8'b11000110; // **   **
            11'h015: data = 8'b11001110; // **  ***
            11'h016: data = 8'b11011110; // ** ****
            11'h017: data = 8'b11110110; // **** **
            11'h018: data = 8'b11100110; // ***  **
            11'h019: data = 8'b11000110; // **   **
            11'h01a: data = 8'b11000110; // **   **
            11'h01b: data = 8'b01111100; //  *****
            11'h01c: data = 8'b00000000; //
            11'h01d: data = 8'b00000000; //
            11'h01e: data = 8'b00000000; //
            11'h01f: data = 8'b00000000; //
            //code x31
            11'h020: data = 8'b00000000; //
            11'h021: data = 8'b00000000; //
            11'h022: data = 8'b00011000; //
            11'h023: data = 8'b00111000; //
            11'h024: data = 8'b01111000; //    **
            11'h025: data = 8'b00011000; //   ***
            11'h026: data = 8'b00011000; //  ****
            11'h027: data = 8'b00011000; //    **
            11'h028: data = 8'b00011000; //    **
            11'h029: data = 8'b00011000; //    **
            11'h02a: data = 8'b00011000; //    **
            11'h02b: data = 8'b01111110; //    **
            11'h02c: data = 8'b00000000; //    **
            11'h02d: data = 8'b00000000; //  ******
            11'h02e: data = 8'b00000000; //
            11'h02f: data = 8'b00000000; //
            //code x32
            11'h030: data = 8'b00000000; //
            11'h031: data = 8'b00000000; //
            11'h032: data = 8'b01111100; //  *****
            11'h033: data = 8'b11000110; // **   **
            11'h034: data = 8'b00000110; //      **
            11'h035: data = 8'b00001100; //     **
            11'h036: data = 8'b00011000; //    **
            11'h037: data = 8'b00110000; //   **
            11'h038: data = 8'b01100000; //  **
            11'h039: data = 8'b11000000; // **
            11'h03a: data = 8'b11000110; // **   **
            11'h03b: data = 8'b11111110; // *******
            11'h03c: data = 8'b00000000; //
            11'h03d: data = 8'b00000000; //
            11'h03e: data = 8'b00000000; //
            11'h03f: data = 8'b00000000; //
            //code x33
            11'h040: data = 8'b00000000; //
            11'h041: data = 8'b00000000; //
            11'h042: data = 8'b01111100; //  *****
            11'h043: data = 8'b11000110; // **   **
            11'h044: data = 8'b00000110; //      **
            11'h045: data = 8'b00000110; //      **
            11'h046: data = 8'b00111100; //   ****
            11'h047: data = 8'b00000110; //      **
            11'h048: data = 8'b00000110; //      **
            11'h049: data = 8'b00000110; //      **
            11'h04a: data = 8'b11000110; // **   **
            11'h04b: data = 8'b01111100; //  *****
            11'h04c: data = 8'b00000000; //
            11'h04d: data = 8'b00000000; //
            11'h04e: data = 8'b00000000; //
            11'h04f: data = 8'b00000000; //
            //code x34
            11'h050: data = 8'b00000000; //
            11'h051: data = 8'b00000000; //
            11'h052: data = 8'b00001100; //     **
            11'h053: data = 8'b00011100; //    ***
            11'h054: data = 8'b00111100; //   ****
            11'h055: data = 8'b01101100; //  ** **
            11'h056: data = 8'b11001100; // **  **
            11'h057: data = 8'b11111110; // *******
            11'h058: data = 8'b00001100; //     **
            11'h059: data = 8'b00001100; //     **
            11'h05a: data = 8'b00001100; //     **
            11'h05b: data = 8'b00011110; //    ****
            11'h05c: data = 8'b00000000; //
            11'h05d: data = 8'b00000000; //
            11'h05e: data = 8'b00000000; //
            11'h05f: data = 8'b00000000; //
            //code x35
            11'h060: data = 8'b00000000; //
            11'h061: data = 8'b00000000; //
            11'h062: data = 8'b11111110; // *******
            11'h063: data = 8'b11000000; // **
            11'h064: data = 8'b11000000; // **
            11'h065: data = 8'b11000000; // **
            11'h066: data = 8'b11111100; // ******
            11'h067: data = 8'b00000110; //      **
            11'h068: data = 8'b00000110; //      **
            11'h069: data = 8'b00000110; //      **
            11'h06a: data = 8'b11000110; // **   **
            11'h06b: data = 8'b01111100; //  *****
            11'h06c: data = 8'b00000000; //
            11'h06d: data = 8'b00000000; //
            11'h06e: data = 8'b00000000; //
            11'h06f: data = 8'b00000000; //
            //code x36
            11'h070: data = 8'b00000000; //
            11'h071: data = 8'b00000000; //
            11'h072: data = 8'b00111000; //   ***
            11'h073: data = 8'b01100000; //  **
            11'h074: data = 8'b11000000; // **
            11'h075: data = 8'b11000000; // **
            11'h076: data = 8'b11111100; // ******
            11'h077: data = 8'b11000110; // **   **
            11'h078: data = 8'b11000110; // **   **
            11'h079: data = 8'b11000110; // **   **
            11'h07a: data = 8'b11000110; // **   **
            11'h07b: data = 8'b01111100; //  *****
            11'h07c: data = 8'b00000000; //
            11'h07d: data = 8'b00000000; //
            11'h07e: data = 8'b00000000; //
            11'h07f: data = 8'b00000000; //
            //code x37
            11'h080: data = 8'b00000000; //
            11'h081: data = 8'b00000000; //
            11'h082: data = 8'b11111110; // *******
            11'h083: data = 8'b11000110; // **   **
            11'h084: data = 8'b00000110; //      **
            11'h085: data = 8'b00000110; //      **
            11'h086: data = 8'b00001100; //     **
            11'h087: data = 8'b00011000; //    **
            11'h088: data = 8'b00110000; //   **
            11'h089: data = 8'b00110000; //   **
            11'h08a: data = 8'b00110000; //   **
            11'h08b: data = 8'b00110000; //   **
            11'h08c: data = 8'b00000000; //
            11'h08d: data = 8'b00000000; //
            11'h08e: data = 8'b00000000; //
            11'h08f: data = 8'b00000000; //
            //code x38
            11'h090: data = 8'b00000000; //
            11'h091: data = 8'b00000000; //
            11'h092: data = 8'b01111100; //  *****
            11'h093: data = 8'b11000110; // **   **
            11'h094: data = 8'b11000110; // **   **
            11'h095: data = 8'b11000110; // **   **
            11'h096: data = 8'b01111100; //  *****
            11'h097: data = 8'b11000110; // **   **
            11'h098: data = 8'b11000110; // **   **
            11'h099: data = 8'b11000110; // **   **
            11'h09a: data = 8'b11000110; // **   **
            11'h09b: data = 8'b01111100; //  *****
            11'h09c: data = 8'b00000000; //
            11'h09d: data = 8'b00000000; //
            11'h09e: data = 8'b00000000; //
            11'h09f: data = 8'b00000000; //
            //code x39
            11'h100: data = 8'b00000000; //
            11'h101: data = 8'b00000000; //
            11'h102: data = 8'b01111100; //  *****
            11'h103: data = 8'b11000110; // **   **
            11'h104: data = 8'b11000110; // **   **
            11'h105: data = 8'b11000110; // **   **
            11'h106: data = 8'b01111110; //  ******
            11'h107: data = 8'b00000110; //      **
            11'h108: data = 8'b00000110; //      **
            11'h109: data = 8'b00000110; //      **
            11'h10a: data = 8'b00001100; //     **
            11'h10b: data = 8'b01111000; //  ****
            11'h10c: data = 8'b00000000; //
            11'h10d: data = 8'b00000000; //
            11'h10e: data = 8'b00000000; //
            11'h10f: data = 8'b00000000; //
            //code x41
            11'h120: data = 8'b00000000; //
            11'h121: data = 8'b00000000; //
            11'h122: data = 8'b00010000; //    *
            11'h123: data = 8'b00111000; //   ***
            11'h124: data = 8'b01101100; //  ** **
            11'h125: data = 8'b11000110; // **   **
            11'h126: data = 8'b11000110; // **   **
            11'h127: data = 8'b11111110; // *******
            11'h128: data = 8'b11000110; // **   **
            11'h129: data = 8'b11000110; // **   **
            11'h12a: data = 8'b11000110; // **   **
            11'h12b: data = 8'b11000110; // **   **
            11'h12c: data = 8'b00000000; //
            11'h12d: data = 8'b00000000; //
            11'h12e: data = 8'b00000000; //
            11'h12f: data = 8'b00000000; //
            //code x42
            11'h130: data = 8'b00000000; //
            11'h131: data = 8'b00000000; //
            11'h132: data = 8'b11111100; // ******
            11'h133: data = 8'b01100110; //  **  **
            11'h134: data = 8'b01100110; //  **  **
            11'h135: data = 8'b01100110; //  **  **
            11'h136: data = 8'b01111100; //  *****
            11'h137: data = 8'b01100110; //  **  **
            11'h138: data = 8'b01100110; //  **  **
            11'h139: data = 8'b01100110; //  **  **
            11'h13a: data = 8'b01100110; //  **  **
            11'h13b: data = 8'b11111100; // ******
            11'h13c: data = 8'b00000000; //
            11'h13d: data = 8'b00000000; //
            11'h13e: data = 8'b00000000; //
            11'h13f: data = 8'b00000000; //
            //code x43
            11'h140: data = 8'b00000000; //
            11'h141: data = 8'b00000000; //
            11'h142: data = 8'b00111100; //   ****
            11'h143: data = 8'b01100110; //  **  **
            11'h144: data = 8'b11000010; // **    *
            11'h145: data = 8'b11000000; // **
            11'h146: data = 8'b11000000; // **
            11'h147: data = 8'b11000000; // **
            11'h148: data = 8'b11000000; // **
            11'h149: data = 8'b11000010; // **    *
            11'h14a: data = 8'b01100110; //  **  **
            11'h14b: data = 8'b00111100; //   ****
            11'h14c: data = 8'b00000000; //
            11'h14d: data = 8'b00000000; //
            11'h14e: data = 8'b00000000; //
            11'h14f: data = 8'b00000000; //
            //code x44
            11'h150: data = 8'b00000000; //
            11'h151: data = 8'b00000000; //
            11'h152: data = 8'b11111000; // *****
            11'h153: data = 8'b01101100; //  ** **
            11'h154: data = 8'b01100110; //  **  **
            11'h155: data = 8'b01100110; //  **  **
            11'h156: data = 8'b01100110; //  **  **
            11'h157: data = 8'b01100110; //  **  **
            11'h158: data = 8'b01100110; //  **  **
            11'h159: data = 8'b01100110; //  **  **
            11'h15a: data = 8'b01101100; //  ** **
            11'h15b: data = 8'b11111000; // *****
            11'h15c: data = 8'b00000000; //
            11'h15d: data = 8'b00000000; //
            11'h15e: data = 8'b00000000; //
            11'h15f: data = 8'b00000000; //
            //code x45
            11'h160: data = 8'b00000000; //
            11'h161: data = 8'b00000000; //
            11'h162: data = 8'b11111110; // *******
            11'h163: data = 8'b01100110; //  **  **
            11'h164: data = 8'b01100010; //  **   *
            11'h165: data = 8'b01101000; //  ** *
            11'h166: data = 8'b01111000; //  ****
            11'h167: data = 8'b01101000; //  ** *
            11'h168: data = 8'b01100000; //  **
            11'h169: data = 8'b01100010; //  **   *
            11'h16a: data = 8'b01100110; //  **  **
            11'h16b: data = 8'b11111110; // *******
            11'h16c: data = 8'b00000000; //
            11'h16d: data = 8'b00000000; //
            11'h16e: data = 8'b00000000; //
            11'h16f: data = 8'b00000000; //
            //code x46
            11'h170: data = 8'b00000000; //
            11'h171: data = 8'b00000000; //
            11'h172: data = 8'b11111110; // *******
            11'h173: data = 8'b01100110; //  **  **
            11'h174: data = 8'b01100010; //  **   *
            11'h175: data = 8'b01101000; //  ** *
            11'h176: data = 8'b01111000; //  ****
            11'h177: data = 8'b01101000; //  ** *
            11'h178: data = 8'b01100000; //  **
            11'h179: data = 8'b01100000; //  **
            11'h17a: data = 8'b01100000; //  **
            11'h17b: data = 8'b11110000; // ****
            11'h17c: data = 8'b00000000; //
            11'h17d: data = 8'b00000000; //
            11'h17e: data = 8'b00000000; //
            11'h17f: data = 8'b00000000; //
            //code x47
            11'h180: data = 8'b00000000; //
            11'h181: data = 8'b00000000; //
            11'h182: data = 8'b00111100; //   ****
            11'h183: data = 8'b01100110; //  **  **
            11'h184: data = 8'b11000010; // **    *
            11'h185: data = 8'b11000000; // **
            11'h186: data = 8'b11000000; // **
            11'h187: data = 8'b11011110; // ** ****
            11'h188: data = 8'b11000110; // **   **
            11'h189: data = 8'b11000110; // **   **
            11'h18a: data = 8'b01100110; //  **  **
            11'h18b: data = 8'b00111010; //   *** *
            11'h18c: data = 8'b00000000; //
            11'h18d: data = 8'b00000000; //
            11'h18e: data = 8'b00000000; //
            11'h18f: data = 8'b00000000; //
        endcase

endmodule
